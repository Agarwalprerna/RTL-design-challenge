module BCD_EX3(input [3:0] BCD , output [3:0] y);
 assign y = BCD + 4'd3;
 endmodule